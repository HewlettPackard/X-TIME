`ifndef MATH_INCLUDE
`define MATH_INCLUDE
function int round_up_div(int a, int b);
    return (a + b - 1) / b;
endfunction
`endif
